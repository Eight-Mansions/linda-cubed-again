pBAV        ��   @  ����Z |@   ��������U |@   ��������P |@   ��������P |    ��������F |@   ��������Z |    ��������i |@   ��������_ |@   ��������P |@   ��������p |@   ��������- |`   ��������d |@   ��������F |@   ��������U |@   ��������Z |@   ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������@7      ���-�   � � � � `@7     ���)�   � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � � K@[        �����  � � � � Z@g        �����  � � � � K@[       �����  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � � @O      ��܀k�  � � � �               ������   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  O      ��܀k�  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � � nC      ��ܪk�  � � � �  `C     ��ܪm�  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �   O        �����  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  @C        ���i�  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � � @C        ������  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � � @C        ��׀k�  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  i ` ``      �����_	  � � � �  i`V VV      �����_	  � � � � i`X LL      �����_	  � � � � i H <<      �����_	 	 � � � � ` \ \\      ��р�P	 
 � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � � @O        ���MS
  � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � � `O        ��؀R  � � � �  ` O       ��؀R  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � � @O H      �����P  � � � � @C <G      ��ր�P  � � � � @7  ;      ��ր�P  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � � A [        �����  � � � � d@g        ����P  � � � � A[       �����  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � � @7      ����-�  � � � � `@7     ����-�  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �   �� 
  ���l�rP� (��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        