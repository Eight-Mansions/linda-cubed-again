pBAV       @� �� )  @  ����F |@   ��������d |@   ��������U |@   ��������A |T   ��������J |@   ��������Z |T   ��������F |`   ��������K |@   ��������P |@   ��������K |@   ��������P |   ��������z |@   ��������K |@   ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������   |    ��������d@C      ������   � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               ��        � � � �               ��        � � � �               �����_    � � � �               ��        � � � �               �����_    � � � �               �����_    � � � � *C        ������  � � � �  KC       ������  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  @[        ����-�  � � � �  @g        ����-�  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � � TO  ;      ������  � � � � sTO <G      ������  � � � � nTO HS      ������  � � � � iTO T      ������  � � � � T O ;      ������  � � � � T O<G      ������  � � � � T OHS      ������  � � � � T OT      ������  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � � `C        ������  � � � �  C       ������  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � � @g O      ������  � � � � @[ CN      ������  � � � � @O  B      ������  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  JC        ����,�  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  @[        ��ڀ��  � � � � 2 [	       ��ڀ��  � � � � 2[       ��ڀ��  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  @O  B    ������  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               ��       � � � �               ��       � � � �               �����_   � � � �               �����_   � � � �               ��       � � � �               ��       � � � � i@O        ������	  � � � � @7        ����+�	  � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �  @O        ������
  � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �  P E EE      ������ 	 � � � �  P`; <<      ������ 
 � � � �  `F FF      ������  � � � �   8 88      ������  � � � �  TR RR      ������  � � � �  d4L @@      ������  � � � �  d@L >>      ������  � � � �  P`D DD      ������ 	 � � � � d@< )0    ��� �_  � � � � d@7 $$    ��� �_  � � � � ZV JJ      �����_  � � � � Z U II      �����_  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  @[        ��ڀ��  � � � �  2 [	       ��ڀ��  � � � �  2[       ��ڀ��  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �   �
"�0�  X B� � � � � p
^���                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  