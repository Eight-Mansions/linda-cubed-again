pBAV       �� ��  	 @  ����_ @   ��������d @   ��������d @   ��������_ @   ��������_ @   ��������_ @   ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������  @< $$      �����_   � � � � p@2 &&      �����_   � � � �  &8 ..      �����_   � � � � F< 11      ����P   � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � � OC ##      ����O  � � � �  <C ''      ����O  � � � �  C **      ����O  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  @        �����O  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � � `C        �����_  � � � �  7        ��� �_  � � � �  @7       ����_  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  `C        �����_  � � � �   C        �����_ 	 � � � �  C       �����_ 	 � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  `C        �����_  � � � �   C        �����_ 	 � � � �  C       �����_ 	 � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �   :NB�bx
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            