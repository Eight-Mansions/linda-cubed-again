pBAV       ��  �� 	  @  ����} @   ��������s @   ��������n @   ��������s @   ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       �������� @7        �� ,�   � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               �����_    � � � �               �����_    � � � �   (C        ��� ��  � � � �   YC       ��� ��  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               �����_   � � � �  x<C        ��� ��  � � � �  xDO        ��� ��  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  @0 $$      ��� ��  � � � �  @2 &&      ��� ��  � � � �  d62 66      ��� ��  � � � �   * **      ��� ��  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �   �4H"��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                