pBAV       @� �� 	  @  ����h �@   ��������h �@   �������� �   ��������M �@   ��������_ �@   ��������H �@   ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    �������� @+        ����LP   � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �  @C        ��ʀ�O  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  [        �����_  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  @+  6      �����_  � � � �  @7 7      �����_  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  @C        �����_  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �   H HH      ������  � � � �  @J JJ      ������  � � � �  L LL      ������  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �   @���\T                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                