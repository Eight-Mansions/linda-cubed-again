pBAV       � ��   @  ���� �@   �������� �@   �������� �@   �������� �@   �������� �@   �������� �@   �������� �@   ��������
 �@   ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������  @+        ��ŀf�   � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �  @C C      ��׀l�  � � � �  @C  B      ��׀l�  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  @C      ��耫�  � � � �  ` C     ��耬�  � � � �  VC     ��耭�  � � � �  n@O      ��耫�  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  @C      ��ـ��  � � � �  ` C
     ��ـ��  � � � �  VC     ��ـ��  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  @C        ��ڀ+�  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  @C      ����k�  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  @O        ������  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �   n`* **      ������  � � � �   `. ..      ������ 	 � � � �  2] QQ      ������ 
 � � � �   d@$ $$      ������  � � � �  d@( ((      ������  � � � �  d E 99      ������  � � � �  d`@ 11      ������  � � � �    ) ))      ������  � � � �   d@- --      ������  � � � �   `0 00      ������  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �   ��*|��r��$�2�@�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              