pBAV        � ��   @  ����M c    ��������M c   ��������W c6   ��������G c@   ��������M c@   ��������W c@   ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������  C :[      ��Հ��   � � � �   7  9      ��Հ��   � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �  C;[      ��Հ��  � � � �  7 :      ��Հ��  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  6O        ����-�  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �   @7        ������ 	 � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  @[ RX      ����  � � � �  @C  E      ����  � � � �  @O IQ      ���� 
 � � � �  @C FH      ����  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �   x@$ $$      ������  � � � �    % %%      ������  � � � �   `& &&      ��� �_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �   ���r��B>,�V                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      