pBAV       �� ��
   @  ���� T@   �������� T@   ��������n TT   ��������< T@   ��������n TT   ��������Z T@   ��������K T@   ��������7 T    ��������f T@   ��������n TT   ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������   T    ��������@[        ��؀)�   � � � �  n [	       ��؀,�   � � � �  @[       ��؀-�   � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � � @O      ��ƀ��  � � � �  T O	     ��ƀ��  � � � �  @O     ��ƀ��  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � � T[        �����  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � � [        ����k�  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � � nTO IQ      ��؀m�  � � � � ZTC <H      ������  � � � � ZTC  ;      ��䀫�  � � � � nTO R      ��䀭�  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � � v[        ����k�  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  @        ��Ȁk�  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  C;[      ��Հ��  � � � �  7 :      ��Հ��  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  Z`* **      ������ 	 � � � � F`? 11      ���n� 
 � � � � <T( ((      ������  � � � �  U@$ $$      ������  � � � � F@& &&      ������  � � � � R*6 66      ������  � � � �  @`7 ++      ������  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � � nTO        ��䀭�	  � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �   (r �8�� ��$����LD"�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             