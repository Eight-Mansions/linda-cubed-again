pBAV       0 ��   @  ����T c    ��������* c   ��������T c@   ��������4 c@   ��������` c@   ��������R c@   ��������R c@   ��������` c@   ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������   c    ��������@O        ��Հ��   � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � � @O O      ��р��  � � � � @C CN      ��р��  � � � � @7  B      ��р��  � � � �               ������   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � � @C        ����f�  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  O        ������  � � � � O       ������  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � � @C      ��؀��  � � � �  ` C	     ��؀��  � � � �  @C     ��؀��  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � � @7        ����  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � � @+        ������ 	 � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � � `T+ ++      ������ 
 � � � � `( ((      ������  � � � � ` ! !!      ������  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �   F 
  �
�	f�	 �`                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      