pBAV       @� ��   @  ����Z �    ��������Z �   ��������f �@   ��������E �    ��������1 �   ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    �������� C <[      ������   � � � �  7 0;      ������   � � � �  +  /      ������   � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � � C ;[      ������  � � � � 7  :      ������  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � � @C  I    ����*�  � � � � @O J    ����*�  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �   C	 I    ����*�  � � � �   O	J    ����*�  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  C I    ����*�  � � � �  OJ    ����*�  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �   ~�����	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                