pBAV       � ��
   @  ����P �T   ��������d �@   ��������P �@   ��������A �@   ��������F �J   ��������K �V   ��������K �    ��������Q �@   ��������Q �@   ��������Z �@   ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������`O T      ����-�   � � � � `C HS      ������   � � � � `C  G      ������   � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �  @        �����P  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � � @+        ��ʀR  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � � @C      ��ڀR  � � � � `@C     ��ڀ.�  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � � HC        ��ր�P  � � � �  ` C       ��ր��  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � � VC        ����R  � � � �  ` C       ����.�  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  O        ����R  � � � �  `O       ����.�  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � � @O        �����_  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � � HC        ��ր�P  � � � �  ` C       ��ր��  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  `@0 $$      �����_	 	 � � � � n@& &&      �����_	 
 � � � � i*$ 00      �����_	 
 � � � � i4$ --      �����_	 
 � � � � iK$ //      �����_	 
 � � � � iT% ++      �����_	 
 � � � � s 6 66      �����_	  � � � � ` **      �����_	 
 � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �   (�� ��2�LL�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      