pBAV         ��
 � F @  ���� @   �������� @   �������� @   �������� @   �������� @   �������� @   �������� @   �������� @   �������� @   �������� @   ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       �������� @< $$      �����_   � � � �   @5 $$      �����_   � � � �  @= %%      �����_   � � � �   @6 %%      �����_   � � � �  @> &&      �����_   � � � �   @7 &&      �����_   � � � �  @? ''      �����_   � � � �   @8 ''      �����_   � � � �  @@ ((      �����_   � � � �   @9 ((      �����_   � � � �  @A ))      �����_   � � � �   @: ))      �����_   � � � �  @B **      �����_   � � � �   @; **      �����_   � � � �  @C ++      �����_   � � � �   @< ++      �����_   � � � �  @< $$      �����_ 	 � � � �   @5 $$      �����_ 	 � � � �  @= %%      �����_ 
 � � � �   @6 %%      �����_ 
 � � � �  @> &&      �����_  � � � �   @7 &&      �����_  � � � �  @? ''      �����_  � � � �   @8 ''      �����_  � � � �  @@ ((      �����_  � � � �   @9 ((      �����_  � � � �  @A ))      �����_  � � � �   @: ))      �����_  � � � �  @B **      �����_  � � � �   @; **      �����_  � � � �               �����_   � � � �               �����_   � � � �  @< $$      �����_  � � � �   @5 $$      �����_  � � � �  @= %%      �����_  � � � �   @6 %%      �����_  � � � �  @> &&      �����_  � � � �   @7 &&      �����_  � � � �  @? ''      �����_  � � � �   @8 ''      �����_  � � � �  @@ ((      �����_  � � � �   @9 ((      �����_  � � � �  @A ))      �����_  � � � �   @: ))      �����_  � � � �  @B **      �����_  � � � �   @; **      �����_  � � � �  @C ++      �����_  � � � �   @< ++      �����_  � � � �  @< $$      �����_  � � � �   @5 $$      �����_  � � � �  @= %%      �����_  � � � �   @6 %%      �����_  � � � �  @> &&      �����_  � � � �   @7 &&      �����_  � � � �  @? ''      �����_  � � � �   @8 ''      �����_  � � � �  @@ ((      �����_  � � � �   @9 ((      �����_  � � � �  @A ))      �����_  � � � �   @: ))      �����_  � � � �  @B **      �����_  � � � �   @; **      �����_  � � � �               �����_   � � � �               �����_   � � � �  @< $$      �����_  � � � �   @5 $$      �����_  � � � �  @= %%      �����_   � � � �   @6 %%      �����_   � � � �  x@> &&      �����_ ! � � � �   @7 &&      �����_ ! � � � �  @? ''      �����_ " � � � �   @8 ''      �����_ " � � � �  @@ ((      �����_ # � � � �   @9 ((      �����_ # � � � �  @A ))      �����_ $ � � � �   @: ))      �����_ $ � � � �  @B **      �����_ % � � � �   @; **      �����_ % � � � �  @C ++      �����_ & � � � �   @< ++      �����_ & � � � �  @< $$      �����_ ' � � � �   @5 $$      �����_ ' � � � �  @= %%      �����_ ( � � � �   @6 %%      �����_ ( � � � �  @> &&      �����_ ) � � � �   @7 &&      �����_ ) � � � �  @? ''      �����_ * � � � �   @8 ''      �����_ * � � � �  @@ ((      �����_ + � � � �   @9 ((      �����_ + � � � �  @A ))      �����_ , � � � �   @: ))      �����_ , � � � �  @B **      �����_ - � � � �   @; **      �����_ - � � � �               �����_   � � � �               �����_   � � � �  @< $$      �����_ . � � � �   @5 $$      �����_ . � � � �  @= %%      �����_ / � � � �   @6 %%      �����_ / � � � �  @> &&      �����_ 0 � � � �   @7 &&      �����_ 0 � � � �  @? ''      �����_ 1 � � � �   @8 ''      �����_ 1 � � � �  @@ ((      �����_ 2 � � � �   @9 ((      �����_ 2 � � � �  @A ))      �����_ 3 � � � �   @: ))      �����_ 3 � � � �  @B **      �����_ 4 � � � �   @; **      �����_ 4 � � � �  @C ++      �����_ 5 � � � �   @< ++      �����_ 5 � � � �  @< $$      �����_ 6 � � � �   @5 $$      �����_ 6 � � � �  @= %%      �����_ 7 � � � �   @6 %%      �����_ 7 � � � �  @> &&      �����_ 8 � � � �   @7 &&      �����_ 8 � � � �  @? ''      �����_ 9 � � � �   @8 ''      �����_ 9 � � � �  @@ ((      �����_ : � � � �   @9 ((      �����_ : � � � �  @A ))      �����_ ; � � � �   @: ))      �����_ ; � � � �  @B **      �����_ < � � � �   @; **      �����_ < � � � �               �����_   � � � �               �����_   � � � �  @< $$      �����_ = � � � �   @5 $$      �����_ = � � � �  @= %%      �����_ > � � � �   @6 %%      �����_ > � � � �  @> &&      �����_ ? � � � �   @7 &&      �����_ ? � � � �  @? ''      �����_ @ � � � �   @8 ''      �����_ @ � � � �  @@ ((      �����_ A � � � �   @9 ((      �����_ A � � � �  @A ))      �����_ B � � � �   @: ))      �����_ B � � � �  @B **      �����_ C � � � �   @; **      �����_ C � � � �  @C ++      �����_ D � � � �   @< ++      �����_ D � � � �  @< $$      �����_	 E � � � �   @5 %%      �����_	 E � � � �  @= &&      �����_	 F � � � �   @6 ''      �����_	 F � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �   ���������������������d*��,"����B$������Pdb�����~���R���������Z����D                                                                                                                                                                                                                                                                                                                                                                                  