pBAV       � ��
   @  ����T �@   ��������@ �   ��������F �6   ��������J �    ��������7 �@   ��������J �@   ��������P �@   ��������2 �@   ��������` �@   �������� �@   ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    ��������   �    �������� JO        ����P   � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �  @C        �����K  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  @C        �����K  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  `@7        ���LL  � � � �  d@C        �����K  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  @O        �����_  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �   @        ���FN  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  @O        ��׀�L  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  @O        �����P  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �   x I II      �����_  � � � �   x L LL      �����_ 	 � � � �   d J JJ      �����_ 
 � � � �   n`G GG      �����_  � � � �   ``H HH      �����_  � � � �   ``V VV      �����_  � � � �   nY YY      �����_  � � � �  s         �����_  � � � �  s       �����_  � � � �  s % %%      �����_  � � � �  i`& &&      �����_  � � � �  n@< 00      �����_  � � � �  n@C <E      �����_  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  @O        ����lN	  � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �   
p�`� &�b�� ^� ��b*�	�(                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      